package axi_test_pkg;

   `include "uvm_macros.svh"
    import uvm_pkg::*;

    import axi_pkg::*;


    `include "axi_write_test.sv"
    `include "axi_read_test.sv"
    `include "axi_MWR_test.sv"

    

endpackage //axi_test_pkg

