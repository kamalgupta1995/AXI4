
package axi_pkg;


import uvm_pkg::*;
`include "uvm_macros.svh"

`define AXI_DATA_WIDTH 256

`include "axi_constants.sv"

`include "axi_config.sv"
`include "bus_enum.sv"
//include files bottom to top
`include "axi_if.sv"
`include "axi_trans.sv"
`include "axi_master_sequencer.sv"
`include "axi_master_driver.sv"
`include "axi_master_monitor.sv"
//`include "axi_slave_driver.sv"
`include "axi_master_agent.sv"
`include "axi_slave_monitor.sv"
`include "axi_slave_agent.sv"
`include "axi_scoreboard.sv"
`include "axi_env.sv"

//`include "axi_seq_lib.sv"
//`include "axi_reset_seq.sv"
`include "axi_Wsequence.sv"
`include "axi_sanity_test.sv"
`include "axi_Rsequence.sv"
`include "axi_read_test.sv"
`include "axi_MWR_sequence.sv"
`include "axi_MWR_test.sv"

`include "axi_tb_top.sv"

endpackage 
